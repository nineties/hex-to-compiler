; plisp2 -- simple lisp interpreter
; Copyright (C) 2026 nineties

(include "std.sv")

; === Memory Allocation

(fun align (n) ; align n to 4-byte boundary
    (return (& (+ n 7) 0xfffffff8))
    )

(def HEAP_BLOCK_SIZE (* 128 (* 1024 1024))) ; 128 MB
(long heap_root)
(long heap_end)
(long heap_pos)
(fun init_heap ()
    (var addr (mmap2 0 HEAP_BLOCK_SIZE
        (| PROT_READ PROT_WRITE)
        (| MAP_PRIVATE MAP_ANONYMOUS)
        -1 0))
    (if (u>= addr 0xfffff001) (do
        (eputs "mmap2 failed\n")
        (exit 1)
        ))
    (= heap_root addr)
    (= heap_pos (align addr))
    (= heap_end (+ addr HEAP_BLOCK_SIZE))
    )

(fun allocate (size)
    (= size (align size))
    (if (>= (+ heap_pos size) heap_end) (do
        (eputs "memory allocation error\n")
        (exit 1)
        ))
    (var addr heap_pos)
    (+= heap_pos size)
    (return addr)
    )

; === Utilities

(fun strndup (from size)
    (var to (allocate (+ size 1)))
    (memcpy to from size)
    (setb to size 0)
    (return to)
    )


; === Nodes

(fun box (val)
    (var cell (allocate 4))
    (set cell 0 val)
    (return cell)
    )
(fun unbox (cell) (get cell))

; last 3 bit of address is used to detect node types
; 000  : int
; 001  : nil
; 010  : cons
; 011  : symbol
; 100  : str
; 101  : lambda
; 110  : macro
; 111  : prim

(def Nint 0)
(def Nnil 1)
(def Ncons 2)
(def Nsymbol 3)
(def Nstr 4)
(def Nlambda 5)
(def Nmacro 6)
(def Nprim 7)

(def nil 1)

(fun fprint_tag (fd tag)
    (if (== tag Nint) (fputs fd "int")
    (if (== tag Nnil) (fputs fd "()")
    (if (== tag Ncons) (fputs fd "cons")
    (if (== tag Nsymbol) (fputs fd "symbol")
    (if (== tag Nstr) (fputs fd "string")
    (if (== tag Nlambda) (fputs fd "lambda")
    (if (== tag Nmacro) (fputs fd "macro")
    (if (== tag Nprim) (fputs fd "prim")
        )))))))))

(fun print_tag (tag) (fprint_tag STDOUT tag))
(fun eprint_tag (tag) (fprint_tag STDERR tag))

(fun tag (node) (return (& 0x7 node)))
(fun untag (node) (return (& 0xfffffff8 node)))
(fun check_tag (t node)
    (if (!= t (tag node)) (do
        (eprint_tag t)
        (eputs " is expected\n")
        (exit 1)
        )))
(fun nset (node pos val) (set (untag node) pos val))
(fun nget (node pos) (get (untag node) pos))

(fun make_int (n) (return (<< n 3)))
(fun to_int (node)
    (check_tag Nint node)
    (return (asr node 3))
    )
(fun make_cons (a b)
    (var cons (allocate 8))
    (set cons 0 a)
    (set cons 1 b)
    (return (| cons Ncons))
    )
(fun length (ls)
    (if (== ls nil) (return 0))
    (check_tag Ncons ls)
    (var n 0)
    (while (!= ls nil) (do
        (+= n 1)
        (= ls (cdr ls))
        ))
    (return n)
    )

(fun cons_p (node) (if (== (tag node) Ncons) (return 1) (return 0)))
(fun car (node)
    (check_tag Ncons node)
    (return (get (untag node) 0))
    )
(fun cdr (node)
    (check_tag Ncons node)
    (return (get (untag node) 1))
    )
(fun caar (node) (return (car (car node))))
(fun cadr (node) (return (car (cdr node))))
(fun cdar (node) (return (cdr (car node))))
(fun cddr (node) (return (cdr (cdr node))))
(fun caaar (node) (return (car (car (car node)))))
(fun caadr (node) (return (car (car (cdr node)))))
(fun cadar (node) (return (car (cdr (car node)))))
(fun caddr (node) (return (car (cdr (cdr node)))))
(fun cdaar (node) (return (cdr (car (car node)))))
(fun cdadr (node) (return (cdr (car (cdr node)))))
(fun cddar (node) (return (cdr (cdr (car node)))))
(fun cdddr (node) (return (cdr (cdr (cdr node)))))

(fun setcar (node v)
    (check_tag Ncons node)
    (nset node 0 v)
    (return nil)
    )
(fun setcdr (node v)
    (check_tag Ncons node)
    (nset node 1 v)
    (return nil)
    )

; interning of symbols
(long symbols 0)    ; { sym, next }

(fun make_symbol (s)
    (var iter symbols)
    (while iter (do
        (var s2 (get iter 0))
        (if (streq (symbol_name s2) s) (return s2))
        (= iter (get iter 1))
        ))
    (var sym (| (allocate 4) Nsymbol))
    (nset sym 0 s)

    (var ent (allocate 8))
    (set ent 0 sym)
    (set ent 1 symbols)
    (= symbols ent)
    (return sym)
    )
(fun symbol_name (s)
    (check_tag Nsymbol s)
    (return (nget s 0))
    )

(long Strue)
(long Sdef)
(long Sset)
(long Sif)
(long Swhile)
(long Sdo)
(long Slambda)
(long Sdefmacro)
(long Squote)
(long Sqquote)
(long Sunquote)
(long Serror)

; variable table
(fun env_push (env sym val)
    (var ent (allocate 12))
    (set ent 0 sym)
    (set ent 1 val)
    (set ent 2 (unbox env))
    (set env ent)
    )

(fun env_update (env sym val)
    (var iter (unbox env))
    (while iter (do
        (if (== (get iter 0) sym) (do
            (set iter 1 val)
            (return)
            ))
        (= iter (get iter 2))
        ))
    (eputs "variable ") (eputs (symbol_name sym)) (eputs " is not found.")
    (exit 1)
    )

(fun env_find (env sym)
    (var iter (unbox env))
    (while iter (do
        (if (== (get iter 0) sym)
            (return (get iter 1)))
        (= iter (get iter 2))
        ))
    (return Serror)
    )

(fun print_env (env)
    (puts "=========\n")
    (var iter (unbox env))
    (while iter (do
        (putx iter) (puts "\n")
        (print_sexp (get iter 0)) (puts " -> ") (print_sexp (get iter 1)) (puts "\n")
        (= iter (get iter 2))
        ))
    (puts "=========\n")
    )

(fun make_quote (e)
    (return (make_cons Squote (make_cons e nil)))
    )
(fun make_qquote (e)
    (return (make_cons Sqquote (make_cons e nil)))
    )
(fun make_unquote (e)
    (return (make_cons Sunquote (make_cons e nil)))
    )


(fun init_symbols ()
    (= Strue (make_symbol "true"))
    (= Sdef (make_symbol "def"))
    (= Sset (make_symbol "set"))
    (= Sif (make_symbol "if"))
    (= Swhile (make_symbol "while"))
    (= Sdo (make_symbol "do"))
    (= Slambda (make_symbol "lambda"))
    (= Sdefmacro (make_symbol "defmacro"))
    (= Squote (make_symbol "quote"))
    (= Sqquote (make_symbol "qquote"))
    (= Sunquote (make_symbol "unquote"))
    (= Serror (make_symbol "error"))
    )

(fun make_str (s)
    (var str (| (allocate 4) Nstr))
    (nset str 0 s)
    (return str)
    )
(fun to_str (s)
    (check_tag Nstr s)
    (return (nget s 0))
    )
(fun make_lambda (env params body)
    (var lam (| (allocate 12) Nlambda))
    (nset lam 0 env)
    (nset lam 1 params)
    (nset lam 2 body)
    (return lam)
    )
(fun make_macro (env params body)
    (var mac (| (allocate 12) Nmacro))
    (nset mac 0 env)
    (nset mac 1 params)
    (nset mac 2 body)
    (return mac)
    )
(fun make_prim (name fun)
    (var prim (| (allocate 8) Nprim))
    (nset prim 0 name)
    (nset prim 1 fun)
    (return prim)
    )

; === Parser and Printer

(fun fprint_str (fd str)
    (fputs fd "\"")
    (while (getb str) (do
        (var c (getb str))
        (var v (escape_char c))
        (if (< v 0)
            (fputc fd c)
            (do
                (fputs fd "\\")
                (fputc fd v)
            ))
        (+= str 1)
        ))
    (fputs fd "\"")
    )

(fun fprint_sexp (fd sexp)
    (var t (tag sexp))
    (if (== t Nint) (fputi fd (to_int sexp))
    (if (== t Nnil) (fputs fd "()")
    (if (== t Ncons) (do
        (fputs fd "(")
        (fprint_sexp fd (car sexp))
        (= sexp (cdr sexp))
        (while (!= sexp nil) (do
            (fputs fd " ")
            (fprint_sexp fd (car sexp))
            (= sexp (cdr sexp))
            ))
        (fputs fd ")")
        )
    (if (== t Nsymbol) (fputs fd (symbol_name sexp))
    (if (== t Nstr) (fprint_str fd (to_str sexp))
    (if (== t Nlambda) (do
        (fputs fd "(lambda ")
        (fprint_sexp fd (nget sexp 0))
        (fputs fd " ...)")
        )
    (if (== t Nmacro) (do
        (fputs fd "(macro ")
        (fprint_sexp fd (nget sexp 0))
        (fputs fd " ...)")
        )
    (if (== t Nprim) (do
        (fputs fd "(prim ")
        (fprint_sexp fd (nget sexp 0))
        (fputs fd " ...)")
        )
        ))))))))
    )
(fun print_sexp (sexp) (fprint_sexp STDOUT sexp))

(fun read_file (path)
    (var fd (open path O_RDONLY))
    (if (< fd 0) (do
        (eputs "open failed: ") (eputs path) (eputs "\n")
        (exit 1)))

    (var file_size (fsize fd))
    (if (< file_size 0) (do
        (eputs "fstat failed: ") (eputs path) (eputs "\n")
        (exit 1)))

    (var buf (allocate (+ file_size 1))) ; +1 for \0
    (var r (read fd buf file_size))
    (if (< r file_size) (do
        (eputs "read failed: ") (eputs path) (eputs "\n")
        (exit 1)
        ))
    (setb buf file_size 0)

    (close fd)
    (return buf)
    )

(fun is_blank (c)
    (if (|| (== c (char " ")) (|| (== c (char "\t")) (== c (char "\n")))) (return 1) (return 0))
    )

(fun skip_spaces_and_comments (textbuf)
    (var addr (unbox textbuf))
    (while (getb addr) (do
        (var c (getb addr))
        (if (== c (char ";"))
            (while (&& (!= (getb addr) (char "\n")) (getb addr)) (+= addr 1))
        (if (is_blank c)
            (+= addr 1)
            (do
                (set textbuf addr)
                (return)
            )))
        ))
    (set textbuf addr)
    )

(fun nextchar (textbuf) (return (getb (unbox textbuf))))

(fun succ (textbuf n)
    (set textbuf (+ (unbox textbuf) n))
    (return textbuf)
    )

(fun is_atom_char (c)
    ; 0-9, a-z, A-Z, +-*/<>=?!_:$%&|^~@[]
    (if (== (getb "xxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxoxxoooxxxooxoxooooooooooooxooooooooooooooooooooooooooooooooxoooxooooooooooooooooooooooooooxoxoxx" c) (char "o"))
        (return 1)
        (return 0)
        )
    )

(fun parse_sym (textbuf)
    (var start (unbox textbuf))
    (while (is_atom_char (nextchar textbuf)) (succ textbuf 1))
    (var end (unbox textbuf))
    (var str (strndup start (- end start)))

    (var c (nextchar textbuf))
    (if (&& (! (is_blank c)) (!= c (char ")"))) (do
        (eputs "junk letters after symbol: ")
        (eputs str)
        (exit 1)
        ))
    (var sym (make_symbol str))
    (return sym)
    )

(fun escape_char (c)
    (if (== c 0) (return (char "0"))
    (if (== c 7) (return (char "a"))
    (if (== c 8) (return (char "b"))
    (if (== c 9) (return (char "t"))
    (if (== c 10) (return (char "n"))
    (if (== c 11) (return (char "v"))
    (if (== c 12) (return (char "f"))
    (if (== c 13) (return (char "r"))
    (if (== c (char "\"")) (return (char "\""))
    (if (== c (char "'")) (return (char "'"))
    (if (== c (char "\\")) (return (char "\\"))
        (return -1)
        ))))))))))))

(fun unescape_char (c)
    (if (== c (char "0")) (return 0)
    (if (== c (char "a")) (return 7)
    (if (== c (char "b")) (return 8)
    (if (== c (char "t")) (return 9)
    (if (== c (char "n")) (return 10)
    (if (== c (char "v")) (return 11)
    (if (== c (char "f")) (return 12)
    (if (== c (char "r")) (return 13)
    (if (== c (char "\"")) (return (char "\"")))
    (if (== c (char "'")) (return (char "'")))
    (if (== c (char "\\")) (return (char "\\"))
        (do
            (eputs "invalid escaped character\n")
            (exit 1)
        )))))))))))

(char[] 4096 parse_str_buf)
(fun parse_str (textbuf)
    (var end parse_str_buf)
    (succ textbuf 1) ; skip '"'
    (while (nextchar textbuf) (do
        (var c (nextchar textbuf))
        (if (== c (char "\"")) (do
            (succ textbuf 1)
            (return (make_str (strndup parse_str_buf (- end parse_str_buf))))
            )
        (if (== c (char "\\")) (do
            (succ textbuf 1)
            (setb end (unescape_char (nextchar textbuf)))
            (+= end 1)
            (succ textbuf 1)
            )
        (do
            (setb end c)
            (+= end 1)
            (succ textbuf 1)
            )))
        ))
    (eputs "invalid string literal: ")
    (eputs parse_str_buf)
    (eputs "\n")
    (exit 1)
    )

(fun parse_uint (textbuf base)
    (var n 0)
    (while (nextchar textbuf) (do
        (var c (nextchar textbuf))
        (var v 0)
        (if (&& (<= (char "0") c) (<= c (char "9")))
            (= v (- c (char "0")))
        (if (&& (<= (char "a") c) (<= c (char "f")))
            (= v (+ (- c (char "a") 10)))
        (if (&& (<= (char "A") c) (<= c (char "F")))
            (= v (+ (- c (char "A") 10)))
            (return (make_int n))
            )))
        (if (>= v base) (do
            (eputs "invalid integer literal\n")
            (exit 1)
            ))
        (= n (+ (* base n) v))
        (succ textbuf 1)
        ))
    (return (make_int n))
    )

(fun parse_int (textbuf)
    (var c (nextchar textbuf))
    (if (! c) (do
        (eputs "invalid integer literal\n")
        (exit 1)
        )
    (if (== c (char "+")) (do
        (succ textbuf 1)
        (return (parse_int textbuf))
        )
    (if (== c (char "-")) (do
        (succ textbuf 1)
        (var v (parse_int textbuf))
        (return (make_int (- (to_int v))))
        )
    (if (== c (char "0")) (do
        (succ textbuf 1)
        (= c (nextchar textbuf))
        (if (== c (char "x"))
            (return (parse_uint (succ textbuf 1) 16))
            )
        (return (parse_uint textbuf 8))
        )))))
    (return (parse_uint textbuf 10))
    )

(fun parse_atom (textbuf)
    (var c (nextchar textbuf))
    (if (== c (char "\""))
        (return (parse_str textbuf))
    (if (&& (>= c (char "0")) (<= c (char "9")))
        (return (parse_int textbuf))
        (return (parse_sym textbuf))
        ))
    )

(fun parse_sexp_list (textbuf)
    (skip_spaces_and_comments textbuf)
    (var c (nextchar textbuf))
    (if (== c 0) (return nil))
    (if (== c (char ")")) (return nil))
    (var sexp (parse_sexp textbuf))
    (var list (parse_sexp_list textbuf))
    (return (make_cons sexp list))
    )

(fun parse_sexp (textbuf)
    (skip_spaces_and_comments textbuf)
    (var addr (unbox textbuf))
    (var c (getb addr))
    (if (== c (char "("))
        (do
            (var ls (parse_sexp_list (succ textbuf 1)))
            (if (!= (nextchar textbuf) (char ")")) (do
                (eputs "syntax error: missing closing parenthesis ')'\n")
                (exit 1)
                ))
            (succ textbuf 1)
            (return ls)
        )
    (if (== c (char "'")) (return (make_quote (parse_sexp (succ textbuf 1))))
    (if (== c (char "`")) (return (make_qquote (parse_sexp (succ textbuf 1))))
    (if (== c (char ",")) (return (make_unquote (parse_sexp (succ textbuf 1))))
        (return (parse_atom textbuf))
        ))))
    )

; === Eval

(fun apply (fn args env)
    (var params (nget fn 0))
    (var body (nget fn 1))
    (var fn_env (box (nget fn 2)))

    ; bind args to params
    (if (== (tag params) Nsymbol)
        (env_push fn_env params args)
        (do
            (if (!= (length params) (length args)) (do
                (eputs "incorrect number of arguments: ")
                (fprint_sexp STDERR params)
                (eputs " <-> ")
                (fprint_sexp STDERR args)
                (eputs "\n")
                (exit 1)
                ))
            (while (!= params nil) (do
                (env_push fn_env (car params) (car args))
                (= params (cdr params))
                (= args (cdr args))
                ))
        ))
    (return (eval_sexp body fn_env))
    )

(fun apply_prim (fn args env)
    (var fp (nget fn 1))
    (var arity (length args))
    (if (== arity 0)
        (return (fp))
    (if (== arity 1)
        (return (fp (car args)))
    (if (== arity 2)
        (return (fp (car args) (cadr args)))
    (if (== arity 3)
        (return (fp (car args) (cadr args) (caddr args)))
        ))))
    (not_implemented "apply_prim")
    )

(fun eval_qquote (sexp env nest)
    (var t (tag sexp))
    (if (!= t Ncons) (return sexp))
    (var head (car sexp))
    (if (== head Squote)
        (return (make_quote (eval_qquote (cadr sexp) env nest)))
    (if (== head Sqquote)
        (return (make_qquote (eval_qquote (cadr sexp) env (+ nest 1))))
    (if (&& (== head Sunquote) (== nest 0))
        (return (eval_sexp (cadr sexp) env))
    (if (== head Sunquote)
        (return (make_unquote (eval_qquote (cadr sexp) env (- nest 1))))
        ))))
    (return (make_cons
        (eval_qquote (car sexp) env nest)
        (eval_qquote (cdr sexp) env nest)
        ))
    )

(fun eval_sexp_list (sexp env)
    (if (== sexp nil) (return nil))
    (return (make_cons
        (eval_sexp (car sexp) env)
        (eval_sexp_list (cdr sexp) env)
        )))

(fun eval_cons (sexp env)
    (var head (car sexp))
    ; special forms
    (if (== head Sdef) (do ; (def x e)
        (if (!= (length sexp) 3) (do
            (eputs "malformed def statement: ")
            (fprint_sexp STDERR sexp)
            (eputs "\n")
            (exit 1)
            ))
        (var x (cadr sexp))
        (var e (caddr sexp))
        (check_tag Nsymbol x)
        (= e (eval_sexp e env))
        (env_push env x e)
        (return nil)
        )
    (if (== head Sset) (not_implemented "eval_cons:set")
    (if (== head Sif) (do
        (if (!= (length sexp) 4) (do
            (eputs "malformed if statement: ")
            (fprint_sexp STDERR sexp)
            (eputs "\n")
            (exit 1)
            ))
        (var cond (cadr sexp))
        (var ifthen (caddr sexp))
        (var ifelse (car (cdddr sexp)))
        (var env_old (unbox env))
        (var ret nil)
        (if (== (eval_sexp cond env) nil)
            (= ret (eval_sexp ifthen env))
            (= ret (eval_sexp ifelse env))
            )
        (set env env_old)
        (return ret)
        )
    (if (== head Swhile) (do
        (if (!= (length sexp) 3) (do
            (eputs "malformed while statement: ")
            (fprint_sexp STDERR sexp)
            (eputs "\n")
            (exit 1)
            ))
        (var cond (cadr sexp))
        (var body (caddr sexp))
        (var env_old (unbox env))
        (while (!= (eval_sexp cond env) nil) (do
            (eval_sexp body env)
            (set env env_old)
            ))
        (return nil)
        )
    (if (== head Sdo) (do
        (var args (cdr sexp))
        (while (!= args nil) (do
            (eval_sexp (car args) env)
            (= args (cdr args))
            ))
        (return nil)
        )
    (if (== head Slambda) (do
        (if (|| (!= (length sexp) 3)
            (&& (!= (tag (cadr sexp)) Ncons) (!= (tag (cadr sexp)) Nsymbol))) (do
            (eputs "malformed lambda expression: ")
            (fprint_sexp STDERR sexp)
            (eputs "\n")
            (exit 1)
            ))
        (var params (cadr sexp))
        (var body (caddr sexp))
        (return (make_lambda params body (unbox env)))
        )
    (if (== head Sdefmacro) (do ; (defmacro f params body)
        (if (|| (!= (length sexp) 4)
            (|| (!= (tag (cadr sexp)) Nsymbol)
            (&& (!= (tag (caddr sexp)) Ncons) (!= (tag (caddr sexp)) Nsymbol)))) (do
            (eputs "malformed defmacro statement: ")
            (fprint_sexp STDERR sexp)
            (eputs "\n")
            (exit 1)
            ))
        (var f (cadr sexp))
        (var params (caddr sexp))
        (var body (car (cdddr sexp)))
        (var mac (make_macro params body (unbox env)))
        (env_push env f mac)
        (return nil)
        )
    (if (== head Squote) (return (cadr sexp))
    (if (== head Sqquote) (not_implemented "eval_cons:qquote")
    (if (== head Sunquote) (not_implemented "eval_cons:unquote")
        ))))))))))
    (var fn (eval_sexp (car sexp) env))
    (var args (eval_sexp_list (cdr sexp) env))
    (var t (tag fn))
    (if (== t Nlambda) (return (apply fn args env))
    (if (== t Nprim) (not_implemented "eval_cons:prim")
        ))
    )

(fun eval_sexp (sexp env)
    (print_sexp sexp) (puts "\n")
    (var t (tag sexp))
    (if (== t Ncons) (return (eval_cons sexp env))
    (if (== t Nsymbol) (do
        (var r (env_find env sexp))
        (puts "====\n")
        (print_sexp r) (puts "\n")
        (print_sexp sexp) (puts "\n")
        (if (== r Serror) (do
            (eputs "undefined variable: ")
            (eputs (symbol_name sexp))
            (eputs "\n")
            (exit 1)
            ))
        (return r)
        )))
    (return sexp)
    )

(fun expand_macro (sexp env nest)
    (var t (tag sexp))
    (if (!= t Ncons) (return sexp))
    (var head (car sexp))
    (if (== head Squote) (return sexp)
    (if (== head Sqquote)
        (return (make_qquote (expand_macro (cadr sexp) env (+ nest 1))))
    (if (== head Sunquote)
        (return (make_unquote (expand_macro (cadr sexp) env (- nest 1))))
        )))
    (if (!= nest 0) (return sexp))
    (if (!= (tag head) Nsymbol) (return sexp))
    (var ent (env_find env head))
    (if (== ent Serror) (return sexp))
    (if (!= (tag ent) Nmacro) (return sexp))
    (return (expand_macro (apply ent (cdr sexp) env)) env nest)
    )

(fun eval_file (path env)
    (var textbuf (box (read_file path)))

    (while 1 (do
        (skip_spaces_and_comments textbuf)
        (if (! (nextchar textbuf)) (return))
        (var sexp (parse_sexp textbuf))
        (= sexp (expand_macro sexp env 0))
        (eval_sexp sexp env)
        ))
    )

; === Primitive Functions
(fun prim_put (s)
    (check_tag Nstr s)
    (puts (to_str s))
    (return nil)
    )

(fun add_prim (name f env)
    (var sym (make_symbol name))
    (var p (make_prim sym f))
    (env_push env sym p)
    )

(fun init_prim (env)
    (add_prim "cons" make_cons env)
    (add_prim "car" car env)
    (add_prim "cdr" cdr env)
    (add_prim "setcar" setcar env)
    (add_prim "setcd" setcdr env)
    (add_prim "print" print_sexp env)
    (add_prim "put" prim_put env)
    )


(fun main (argc argv)
    (if (<= argc 1) (do
        (puts "no input file")
        (exit 1)
        ))

    (init_heap)

    (var env (box 0))

    (init_symbols)
    (init_prim env)

    (eval_file "plisp/init.lisp" env)
    (eval_file (get argv 1) env)
    )
