; hello.sv

(include "std.sv")

(fun main ()
    (puts "Hello World!")
    )
